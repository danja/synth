.title KiCad schematic
U1 Net-_R6-Pad2_ Net-_R6-Pad2_ Net-_Q1-Pad1_ NC_01 GND Net-_R5-Pad2_ Net-_R5-Pad2_ Net-_MES1-Pad2_ Net-_R5-Pad1_ Net-_R6-Pad1_ NC_02 Net-_R1-Pad1_ Net-_Q2-Pad1_ Net-_Q2-Pad2_ TL084
R8 Net-_R6-Pad1_ GND 22k
R6 Net-_R6-Pad1_ Net-_R6-Pad2_ 2k2
R5 Net-_R5-Pad1_ Net-_R5-Pad2_ 2k2
R7 Net-_MES1-Pad2_ Net-_R5-Pad1_ 22k
Q1 Net-_Q1-Pad1_ GND +12V 2N3904
Q2 Net-_Q2-Pad1_ Net-_Q2-Pad2_ Net-_Q2-Pad3_ 2N3904
R4 Net-_Q1-Pad1_ Net-_Q2-Pad3_ 10k
R2 Net-_R1-Pad1_ GND 10k
R3 Net-_Q2-Pad1_ -12V 56k
MES1 GND Net-_MES1-Pad2_ Voltmeter_DC
R1 Net-_R1-Pad1_ -12V 10k
.end
